* Created by KLayout

* cell TOP
* pin TP1
* pin Vin2,Vout4
* pin TP2
* pin Vout
* pin VM
* pin VDD
* pin SUBSTRATE
.SUBCKT TOP 7 8 9 11 12 14 16
* net 7 TP1
* net 8 Vin2,Vout4
* net 9 TP2
* net 11 Vout
* net 12 VM
* net 14 VDD
* net 16 SUBSTRATE
* device instance $1 r0 *1 87,73.5 PMOS
M$1 11 10 14 14 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $2 r0 *1 39,73.5 PMOS
M$2 9 7 14 14 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $3 r0 *1 2,73.5 PMOS
M$3 4 4 14 14 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $4 r0 *1 66.5,73.5 PMOS
M$4 15 2 14 14 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $5 r0 *1 19,73.5 PMOS
M$5 7 7 14 14 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $6 r0 *1 28,68.5 PMOS
M$6 8 6 14 14 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $7 r0 *1 8,68.5 PMOS
M$7 6 6 14 14 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $8 r0 *1 75,67.5 PMOS
M$8 10 8 15 14 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $9 r0 *1 59,67.5 PMOS
M$9 2 9 15 14 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $10 r0 *1 75,55 NMOS
M$10 3 8 10 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $11 r0 *1 59,55 NMOS
M$11 3 9 2 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $12 r0 *1 50,55 NMOS
M$12 1 9 9 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $13 r0 *1 33.5,55 NMOS
M$13 1 9 8 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $14 r0 *1 28,55 NMOS
M$14 1 8 8 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $15 r0 *1 85,55 NMOS
M$15 16 10 11 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $16 r0 *1 44.5,55 NMOS
M$16 1 8 9 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $17 r0 *1 19,55 NMOS
M$17 5 13 7 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $18 r0 *1 8,55 NMOS
M$18 5 12 6 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $19 r0 *1 2,51 NMOS
M$19 16 4 4 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $20 r0 *1 13.5,51 NMOS
M$20 16 4 5 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $21 r0 *1 66.5,47 NMOS
M$21 16 2 3 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $22 r0 *1 39,45.5 NMOS
M$22 16 1 1 16 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
