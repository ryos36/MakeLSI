* Created by KLayout

* cell TOP
* pin VM
* pin VSS
.SUBCKT TOP 3 4
* net 3 VM
* net 4 VSS
* device instance $1 r0 *1 8,55 NMOS
M$1 4 3 2 4 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $2 r0 *1 2,51 NMOS
M$2 4 1 1 4 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
