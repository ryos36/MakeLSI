.title KiCad schematic
M1 Net-_M1-Pad1_ Net-_M1-Pad1_ /VDD /VDD PMOS l=1u w=2u
M2 Net-_M1-Pad1_ Net-_M1-Pad1_ /VSS /VSS NMOS l=1u w=2u
M3 Net-_M3-Pad1_ /VM Net-_M3-Pad3_ /VSS NMOS l=1u w=2u
M4 Net-_M3-Pad1_ Net-_M3-Pad1_ /VDD /VDD PMOS l=1u w=2u
M5 Net-_M3-Pad3_ Net-_M1-Pad1_ /VSS /VSS NMOS l=1u w=2u
M6 Net-_M12-Pad2_ Net-_M12-Pad2_ /VDD /VDD PMOS l=1u w=2u
M7 Net-_M12-Pad2_ /VP Net-_M3-Pad3_ /VSS NMOS l=1u w=2u
M8 Net-_M11-Pad1_ Net-_M3-Pad1_ /VDD /VDD PMOS l=1u w=2u
*M9 Net-_M11-Pad1_ Net-_M11-Pad1_ Net-_M10-Pad1_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M20 Net-_M19-Pad1_ Net-_M11-Pad1_ Net-_M16-Pad3_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M18 Net-_M16-Pad3_ Net-_M15-Pad1_ Net-_M10-Pad3_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M16 Net-_M15-Pad1_ Net-_M11-Pad2_ Net-_M16-Pad3_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M22 /Vout Net-_M19-Pad1_ Net-_M10-Pad3_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M11 Net-_M11-Pad1_ Net-_M11-Pad2_ Net-_M10-Pad1_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M10 Net-_M10-Pad1_ Net-_M10-Pad1_ Net-_M10-Pad3_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M13 Net-_M11-Pad2_ Net-_M11-Pad1_ Net-_M10-Pad1_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M14 Net-_M11-Pad2_ Net-_M11-Pad2_ Net-_M10-Pad1_ Net-_M10-Pad3_ NMOS l=1u w=2u
*M19 Net-_M19-Pad1_ Net-_M11-Pad1_ Net-_M15-Pad3_ /VDD PMOS l=1u w=6u
*M17 Net-_M15-Pad3_ Net-_M15-Pad1_ /VDD /VDD PMOS l=1u w=2u
*M15 Net-_M15-Pad1_ Net-_M11-Pad2_ Net-_M15-Pad3_ /VDD PMOS l=1u w=2u
*M21 /Vout Net-_M19-Pad1_ /VDD /VDD PMOS l=1u w=17u
*M12 Net-_M11-Pad2_ Net-_M12-Pad2_ /VDD /VDD PMOS l=1u w=2u
.end
