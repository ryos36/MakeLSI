*

.subckt cc_osc


M35 NC-M35-0 NC-M35-1 NC-M35-2 NC-M35-3 PMOS_OR1 l=1u w=6u
M34 NC-M34-0 NC-M34-1 NC-M34-2 NC-M34-3 NMOS_OR1 l=1u w=2u
M32 NC-M32-0 NC-M32-1 NC-M32-2 NC-M32-3 PMOS_OR1 l=1u w=6u
M33 NC-M33-0 NC-M33-1 NC-M33-2 NC-M33-3 NMOS_OR1 l=1u w=2u
M27 NC-M27-0 NC-M27-1 NC-M27-2 NC-M27-3 NMOS_OR1 l=1u w=2u
M37 NC-M37-0 NC-M37-1 NC-M37-2 NC-M37-3 PMOS_OR1 l=1u w=6u
M36 NC-M36-0 NC-M36-1 NC-M36-2 NC-M36-3 NMOS_OR1 l=1u w=2u
M31 NC-M31-0 NC-M31-1 NC-M31-2 NC-M31-3 NMOS_OR1 l=1u w=2u
M28 NC-M28-0 NC-M28-1 NC-M28-2 NC-M28-3 NMOS_OR1 l=1u w=2u
M30 NC-M30-0 NC-M30-1 NC-M30-2 NC-M30-3 PMOS_OR1 l=1u w=6u
M29 NC-M29-0 NC-M29-1 NC-M29-2 NC-M29-3 NMOS_OR1 l=1u w=2u
M49 NC-M49-0 NC-M49-1 NC-M49-2 NC-M49-3 NMOS_OR1 l=1u w=2u
M52 NC-M52-0 NC-M52-1 NC-M52-2 NC-M52-3 PMOS_OR1 l=1u w=6u
M50 NC-M50-0 NC-M50-1 NC-M50-2 NC-M50-3 PMOS_OR1 l=1u w=6u
M48 NC-M48-0 NC-M48-1 NC-M48-2 NC-M48-3 NMOS_OR1 l=1u w=2u
M51 NC-M51-0 NC-M51-1 NC-M51-2 NC-M51-3 NMOS_OR1 l=1u w=2u
M42 NC-M42-0 NC-M42-1 NC-M42-2 NC-M42-3 PMOS_OR1 l=1u w=6u
M40 NC-M40-0 NC-M40-1 NC-M40-2 NC-M40-3 PMOS_OR1 l=1u w=6u
M38 NC-M38-0 NC-M38-1 NC-M38-2 NC-M38-3 NMOS_OR1 l=1u w=2u
M41 NC-M41-0 NC-M41-1 NC-M41-2 NC-M41-3 NMOS_OR1 l=1u w=2u
M39 NC-M39-0 NC-M39-1 NC-M39-2 NC-M39-3 NMOS_OR1 l=1u w=2u
M43 NC-M43-0 NC-M43-1 NC-M43-2 NC-M43-3 NMOS_OR1 l=1u w=2u
M46 NC-M46-0 NC-M46-1 NC-M46-2 NC-M46-3 NMOS_OR1 l=1u w=2u
M47 NC-M47-0 NC-M47-1 NC-M47-2 NC-M47-3 PMOS_OR1 l=1u w=6u
M44 NC-M44-0 NC-M44-1 NC-M44-2 NC-M44-3 NMOS_OR1 l=1u w=2u
M45 NC-M45-0 NC-M45-1 NC-M45-2 NC-M45-3 PMOS_OR1 l=1u w=6u

.ends
