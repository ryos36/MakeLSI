* Created by KLayout

* cell TOP
* pin OUT
* pin VDD
* pin VSS
.SUBCKT TOP 1 2 3
* net 1 OUT
* net 2 VDD
* net 3 VSS
* device instance $1 r0 *1 -4,0.5 PMOS
M$1 2 1 1 2 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $2 r0 *1 -4,-11 NMOS
M$2 3 1 1 3 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
