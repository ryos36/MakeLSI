* Created by KLayout

* cell TOP
* pin Vin2,Vout2
* pin Vin1,Vout1
* pin Vout4
* pin Vout3
* pin VM
* pin VDD
* pin VSS
.SUBCKT TOP 4 5 6 7 8 10 11
* net 4 Vin2,Vout2
* net 5 Vin1,Vout1
* net 6 Vout4
* net 7 Vout3
* net 8 VM
* net 10 VDD
* net 11 VSS
* device instance $1 r0 *1 39,73.5 PMOS
M$1 7 5 10 10 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $2 r0 *1 2,73.5 PMOS
M$2 2 2 10 10 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $3 r0 *1 19,73.5 PMOS
M$3 5 5 10 10 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $4 r0 *1 28,68.5 PMOS
M$4 6 4 10 10 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $5 r0 *1 8,68.5 PMOS
M$5 4 4 10 10 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $6 r0 *1 50,55 NMOS
M$6 1 7 7 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $7 r0 *1 33.5,55 NMOS
M$7 1 7 6 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $8 r0 *1 28,55 NMOS
M$8 1 6 6 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $9 r0 *1 44.5,55 NMOS
M$9 1 6 7 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $10 r0 *1 19,55 NMOS
M$10 3 9 5 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $11 r0 *1 8,55 NMOS
M$11 3 8 4 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $12 r0 *1 13.5,51 NMOS
M$12 11 2 3 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $13 r0 *1 2,51 NMOS
M$13 11 2 2 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $14 r0 *1 39,45.5 NMOS
M$14 11 1 1 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
