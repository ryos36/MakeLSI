*

.subckt Top
+       FB ; input
+       IN ; input
+       VDD ; input
+       VSS ; input


M2 IN IN VSS VSS NMOS l=1u w=2u
M27 IN IN VSS VSS NMOS l=1u w=2u
M1 IN IN VDD VDD PMOS l=1u w=6u
M3 IN IN VDD VDD PMOS l=1u w=6u
M4 IN FB IN VSS NMOS l=1u w=2u

.ends
