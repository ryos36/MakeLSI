* Created by KLayout

* cell TOP
* pin Vout2
* pin Vout1
* pin Vout
* pin VM
* pin Vin2
* pin Vin1
* pin VDD
* pin VSS
.SUBCKT TOP 9 10 12 13 15 16 17 19
* net 9 Vout2
* net 10 Vout1
* net 12 Vout
* net 13 VM
* net 15 Vin2
* net 16 Vin1
* net 17 VDD
* net 19 VSS
* device instance $1 r0 *1 89.75,73.5 PMOS
M$1 12 11 17 17 PMOS L=1U W=5.5U AS=13.75P AD=13.75P PS=16U PD=16U
* device instance $2 r0 *1 69.5,73.5 PMOS
M$2 18 3 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $3 r0 *1 39,73.5 PMOS
M$3 10 8 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $4 r0 *1 2,73.5 PMOS
M$4 5 5 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $5 r0 *1 19,73.5 PMOS
M$5 8 8 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $6 r0 *1 28,68.5 PMOS
M$6 9 7 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $7 r0 *1 8,68.5 PMOS
M$7 7 7 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $8 r0 *1 78,67.5 PMOS
M$8 11 15 18 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $9 r0 *1 62,67.5 PMOS
M$9 3 16 18 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $10 r0 *1 78,55 NMOS
M$10 4 15 11 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $11 r0 *1 62,55 NMOS
M$11 4 16 3 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $12 r0 *1 50,55 NMOS
M$12 2 10 10 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $13 r0 *1 33.5,55 NMOS
M$13 2 10 9 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $14 r0 *1 88,55 NMOS
M$14 19 11 12 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $15 r0 *1 28,55 NMOS
M$15 2 9 9 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $16 r0 *1 13.5,51 NMOS
M$16 1 5 6 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $17 r0 *1 2,51 NMOS
M$17 19 5 5 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $18 r0 *1 44.5,55 NMOS
M$18 2 9 10 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $19 r0 *1 19,55 NMOS
M$19 6 14 8 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $20 r0 *1 8,55 NMOS
M$20 6 13 7 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $21 r0 *1 69.5,47 NMOS
M$21 19 3 4 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $22 r0 *1 39,45.5 NMOS
M$22 19 2 2 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
