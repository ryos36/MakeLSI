*.TITLE KICAD SCHEMATIC
M1 /X /A /VDD /VDD PMOS L=1U W=6U
M2 /X /A /VSS /VSS NMOS L=1U W=2U
.ENDS
