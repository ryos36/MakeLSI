* Created by KLayout

* cell TOP
* pin IN
* pin OUT
* pin Vin2
* pin VDD
* pin VSS
.SUBCKT TOP 1 21 22 23 25
* net 1 IN
* net 21 OUT
* net 22 Vin2
* net 23 VDD
* net 25 VSS
* device instance $1 r0 *1 -2,18 PMOS
M$1 23 14 14 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $2 r0 *1 19,18 PMOS
M$2 23 16 16 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $3 r0 *1 39,18 PMOS
M$3 23 11 11 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $4 r0 *1 59,18 PMOS
M$4 23 17 17 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $5 r0 *1 79.5,18 PMOS
M$5 23 18 18 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $6 r0 *1 102.5,21.5 PMOS
M$6 7 9 24 23 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $7 r0 *1 118.5,21.5 PMOS
M$7 19 22 24 23 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $8 r0 *1 -1.5,27 PMOS
M$8 23 14 15 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $9 r0 *1 19.5,27 PMOS
M$9 23 16 10 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $10 r0 *1 39.5,27 PMOS
M$10 23 11 12 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $11 r0 *1 59.5,27 PMOS
M$11 23 17 13 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $12 r0 *1 80,27 PMOS
M$12 23 18 9 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $13 r0 *1 110,27.5 PMOS
M$13 24 7 23 23 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $14 r0 *1 130.5,27.5 PMOS
M$14 20 19 23 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $15 r0 *1 146.5,27.5 PMOS
M$15 21 20 23 23 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $16 r0 *1 -12,-4 NMOS
M$16 25 1 1 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $17 r0 *1 -4,-4 NMOS
M$17 25 1 2 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $18 r0 *1 17,-4 NMOS
M$18 25 1 3 25 NMOS L=1U W=2U AS=4P AD=6P PS=8U PD=10U
* device instance $19 r0 *1 37,-4 NMOS
M$19 25 1 4 25 NMOS L=1U W=2U AS=4P AD=6P PS=8U PD=10U
* device instance $20 r0 *1 57,-4 NMOS
M$20 25 1 5 25 NMOS L=1U W=2U AS=4P AD=6P PS=8U PD=10U
* device instance $21 r0 *1 77.5,-4 NMOS
M$21 25 1 6 25 NMOS L=1U W=2U AS=4P AD=6P PS=8U PD=10U
* device instance $22 r0 *1 110,-1 NMOS
M$22 25 7 8 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $23 r0 *1 17,5.5 NMOS
M$23 3 14 16 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $24 r0 *1 23,5.5 NMOS
M$24 3 15 10 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $25 r0 *1 43,5.5 NMOS
M$25 4 10 12 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $26 r0 *1 57,5.5 NMOS
M$26 5 11 17 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $27 r0 *1 83.5,5.5 NMOS
M$27 6 13 9 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $28 r0 *1 102.5,7 NMOS
M$28 8 9 7 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $29 r0 *1 118.5,7 NMOS
M$29 8 22 19 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $30 r0 *1 128.5,7 NMOS
M$30 25 19 20 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $31 r0 *1 144.5,7 NMOS
M$31 25 20 21 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $32 r0 *1 -4,5.5 NMOS
M$32 2 18 14 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $33 r0 *1 2.5,5.5 NMOS
M$33 2 9 15 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $34 r0 *1 37,5.5 NMOS
M$34 4 16 11 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $35 r0 *1 63,5.5 NMOS
M$35 5 12 13 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $36 r0 *1 77.5,5.5 NMOS
M$36 6 17 18 25 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
