* Created by KLayout

* cell TOP
* pin IN
* pin OUT
* pin Vin2
* pin VDD
* pin VSS
.SUBCKT TOP 1 20 21 22 24
* net 1 IN
* net 20 OUT
* net 21 Vin2
* net 22 VDD
* net 24 VSS
* device instance $1 r0 *1 -2,18 PMOS
M$1 22 14 14 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $2 r0 *1 19,18 PMOS
M$2 22 16 16 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $3 r0 *1 39,18 PMOS
M$3 22 11 11 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $4 r0 *1 59,18 PMOS
M$4 22 17 17 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $5 r0 *1 79.5,18 PMOS
M$5 22 18 18 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $6 r0 *1 102.5,21.5 PMOS
M$6 7 9 23 22 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $7 r0 *1 118.5,21.5 PMOS
M$7 19 21 23 22 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $8 r0 *1 -1.5,27 PMOS
M$8 22 14 15 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $9 r0 *1 19.5,27 PMOS
M$9 22 16 10 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $10 r0 *1 39.5,27 PMOS
M$10 22 11 12 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $11 r0 *1 59.5,27 PMOS
M$11 22 17 13 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $12 r0 *1 80,27 PMOS
M$12 22 18 9 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $13 r0 *1 110,27.5 PMOS
M$13 23 7 22 22 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $14 r0 *1 130.5,27.5 PMOS
M$14 20 19 22 22 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $15 r0 *1 128.5,7 NMOS
M$15 24 19 20 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $16 r0 *1 118.5,7 NMOS
M$16 8 21 19 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $17 r0 *1 102.5,7 NMOS
M$17 8 9 7 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $18 r0 *1 77.5,5.5 NMOS
M$18 6 17 18 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $19 r0 *1 57,5.5 NMOS
M$19 5 11 17 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $20 r0 *1 -12,-4 NMOS
M$20 24 1 1 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $21 r0 *1 -4,-4 NMOS
M$21 24 1 2 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $22 r0 *1 37,-4 NMOS
M$22 24 1 4 24 NMOS L=1U W=2U AS=4P AD=6P PS=8U PD=10U
* device instance $23 r0 *1 17,-4 NMOS
M$23 24 1 3 24 NMOS L=1U W=2U AS=4P AD=6P PS=8U PD=10U
* device instance $24 r0 *1 77.5,-4 NMOS
M$24 24 1 6 24 NMOS L=1U W=2U AS=4P AD=6P PS=8U PD=10U
* device instance $25 r0 *1 63,5.5 NMOS
M$25 5 12 13 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $26 r0 *1 23,5.5 NMOS
M$26 3 15 10 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $27 r0 *1 110,-1 NMOS
M$27 24 7 8 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $28 r0 *1 17,5.5 NMOS
M$28 3 14 16 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $29 r0 *1 83.5,5.5 NMOS
M$29 6 13 9 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $30 r0 *1 57,-4 NMOS
M$30 24 1 5 24 NMOS L=1U W=2U AS=4P AD=6P PS=8U PD=10U
* device instance $31 r0 *1 -4,5.5 NMOS
M$31 2 18 14 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $32 r0 *1 2.5,5.5 NMOS
M$32 2 9 15 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $33 r0 *1 37,5.5 NMOS
M$33 4 16 11 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $34 r0 *1 43,5.5 NMOS
M$34 4 10 12 24 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
