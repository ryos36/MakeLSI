* Created by KLayout

* cell TOP
* pin OUT
* pin VDD
* pin VSS
.SUBCKT TOP 7 8 9
* net 7 OUT
* net 8 VDD
* net 9 VSS
* device instance $1 r0 *1 33.5,0.5 PMOS
M$1 8 5 6 8 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $2 r0 *1 18.5,0.5 PMOS
M$2 8 3 4 8 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $3 r0 *1 41,0.5 PMOS
M$3 8 6 7 8 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $4 r0 *1 11,0.5 PMOS
M$4 8 2 3 8 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $5 r0 *1 26,0.5 PMOS
M$5 8 4 5 8 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $6 r0 *1 3.5,0.5 PMOS
M$6 8 1 2 8 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $7 r0 *1 -4,0.5 PMOS
M$7 8 7 1 8 PMOS L=1U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $8 r0 *1 33.5,-11 NMOS
M$8 9 5 6 9 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $9 r0 *1 26,-11 NMOS
M$9 9 4 5 9 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $10 r0 *1 18.5,-11 NMOS
M$10 9 3 4 9 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $11 r0 *1 41,-11 NMOS
M$11 9 6 7 9 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $12 r0 *1 11,-11 NMOS
M$12 9 2 3 9 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $13 r0 *1 3.5,-11 NMOS
M$13 9 1 2 9 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $14 r0 *1 -4,-11 NMOS
M$14 9 7 1 9 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
