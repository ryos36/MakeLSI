* Created by KLayout

* cell TOP
* pin Vm
* pin Vp
* pin VDD
* pin VSS
.SUBCKT TOP 13 14 17 19
* net 13 Vm
* net 14 Vp
* net 17 VDD
* net 19 VSS
* device instance $1 r0 *1 98,73.5 PMOS
M$1 12 11 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $2 r0 *1 48,73.5 PMOS
M$2 9 7 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $3 r0 *1 2,73.5 PMOS
M$3 1 1 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $4 r0 *1 25,73.5 PMOS
M$4 7 7 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $5 r0 *1 86,68.5 PMOS
M$5 11 8 18 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $6 r0 *1 78.5,73.5 PMOS
M$6 18 3 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $7 r0 *1 71,68.5 PMOS
M$7 3 9 18 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $8 r0 *1 37,68.5 PMOS
M$8 8 6 17 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $9 r0 *1 14,68.5 PMOS
M$9 6 6 16 17 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $10 r0 *1 98,57 NMOS
M$10 19 11 12 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $11 r0 *1 86,57 NMOS
M$11 4 8 11 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $12 r0 *1 37,57 NMOS
M$12 2 8 8 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $13 r0 *1 14,55 NMOS
M$13 5 13 6 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $14 r0 *1 25,55 NMOS
M$14 5 14 7 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $15 r0 *1 19.5,51 NMOS
M$15 19 1 5 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $16 r0 *1 71,57 NMOS
M$16 4 15 3 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $17 r0 *1 2,51 NMOS
M$17 19 1 1 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $18 r0 *1 59,57 NMOS
M$18 2 10 10 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $19 r0 *1 53.5,57 NMOS
M$19 2 8 9 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $20 r0 *1 78.5,49 NMOS
M$20 19 3 4 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $21 r0 *1 42.5,57 NMOS
M$21 2 9 8 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $22 r0 *1 48,49 NMOS
M$22 19 2 2 19 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
