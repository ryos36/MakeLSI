*

.subckt build-vco
+       FB ; input
+       IN ; input
+       OUT ; output
+       VDD ; input
+       VSS ; input


M2 Net-_M2-D_ IN VSS VSS NMOS_OR1 l=1u w=2u
M27 IN IN VSS VSS NMOS_OR1 l=1u w=2u
M1 OUT OUT VDD VDD PMOS_OR1 l=1u w=6u
M3 OUT OUT VDD VDD PMOS_OR1 l=1u w=6u
M4 OUT FB Net-_M2-D_ VSS NMOS_OR1 l=1u w=2u
M5 OUT FB Net-_M2-D_ VSS NMOS_OR1 l=1u w=2u

.ends
