* Created by KLayout

* cell TOP
* pin VDD,VP
* pin VM
* pin VSS
.SUBCKT TOP 1 9 11
* net 1 VDD,VP
* net 9 VM
* net 11 VSS
* device instance $1 r0 *1 39,73.5 PMOS
M$1 7 2 1 1 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $2 r0 *1 2,73.5 PMOS
M$2 5 5 1 1 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $3 r0 *1 19,73.5 PMOS
M$3 2 2 1 1 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $4 r0 *1 28,68.5 PMOS
M$4 3 6 1 1 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $5 r0 *1 8,68.5 PMOS
M$5 6 6 1 1 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $6 r0 *1 33.5,55 NMOS
M$6 4 7 3 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $7 r0 *1 28,55 NMOS
M$7 4 3 3 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $8 r0 *1 19,55 NMOS
M$8 8 10 2 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $9 r0 *1 8,55 NMOS
M$9 8 9 6 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $10 r0 *1 13.5,51 NMOS
M$10 11 5 8 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $11 r0 *1 2,51 NMOS
M$11 11 5 5 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $12 r0 *1 39,47 NMOS
M$12 11 4 4 11 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
