*

.subckt Top
+       IN ; input
+       VDD ; input
+       VSS ; input


M1 IN IN VDD VDD PMOS l=1u w=6u
M27 IN IN VSS VSS NMOS l=1u w=2u

.ends
