*

.subckt build-vco
+       IN ; input
+       VDD ; input
+       VSS ; input


M27 IN IN VSS VSS NMOS_OR1 l=1u w=2u
M1 IN IN VDD VDD PMOS_OR1 l=1u w=6u

.ends
