*

.subckt Top
+       FB ; input
+       IN ; input
+       OUT ; output
+       VDD ; input
+       VSS ; input


M11 Net-_M10-S_ IN VSS VSS NMOS l=1u w=2u
M7 Net-_M10-S_ IN VSS VSS NMOS l=1u w=2u
M4 Net-_M1-D_ FB IN VSS NMOS l=1u w=2u
M3 Net-_M10-G_ Net-_M1-D_ VDD VDD PMOS l=1u w=6u
M5 Net-_M10-G_ OUT IN VSS NMOS l=1u w=2u
M1 Net-_M1-D_ Net-_M1-D_ VDD VDD PMOS l=1u w=6u
M10 Net-_M10-D_ Net-_M10-G_ Net-_M10-S_ VSS NMOS l=1u w=2u
M9 Net-_M10-D_ Net-_M6-D_ VDD VDD PMOS l=1u w=6u
M8 Net-_M6-D_ Net-_M6-D_ VDD VDD PMOS l=1u w=6u
M6 Net-_M6-D_ Net-_M1-D_ Net-_M10-S_ VSS NMOS l=1u w=2u
M27 IN IN VSS VSS NMOS l=1u w=2u
M2 IN IN VSS VSS NMOS l=1u w=2u

.ends
