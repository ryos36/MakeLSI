* Created by KLayout

* cell TOP
* pin VDD,VP
* pin Vout1
* pin Vout2
* pin Vin2
* pin Vin1
* pin VSS
.SUBCKT TOP 1 2 4 5 6 7
* net 1 VDD,VP
* net 2 Vout1
* net 4 Vout2
* net 5 Vin2
* net 6 Vin1
* net 7 VSS
* device instance $1 r0 *1 39,73.5 PMOS
M$1 2 6 1 1 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $2 r0 *1 28,68.5 PMOS
M$2 4 5 1 1 PMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $3 r0 *1 50,55 NMOS
M$3 3 2 2 7 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $4 r0 *1 44.5,55 NMOS
M$4 3 4 2 7 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $5 r0 *1 33.5,55 NMOS
M$5 3 2 4 7 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $6 r0 *1 28,55 NMOS
M$6 3 4 4 7 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
* device instance $7 r0 *1 39,45.5 NMOS
M$7 7 3 3 7 NMOS L=1U W=2U AS=5P AD=5P PS=9U PD=9U
.ENDS TOP
