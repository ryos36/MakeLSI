*

.subckt tb_VCO_buf


M7 NC-M7-0 NC-M7-1 NC-M7-2 NC-M7-3 PMOS_OR1 l=1u w=6u
M5 NC-M5-0 NC-M5-1 NC-M5-2 NC-M5-3 PMOS_OR1 l=1u w=2u
M8 NC-M8-0 NC-M8-1 NC-M8-2 NC-M8-3 NMOS_OR1 l=1u w=2u
M1 NC-M1-0 NC-M1-1 NC-M1-2 NC-M1-3 PMOS_OR1 l=1u w=2u
M3 NC-M3-0 NC-M3-1 NC-M3-2 NC-M3-3 PMOS_OR1 l=1u w=2u
M2 NC-M2-0 NC-M2-1 NC-M2-2 NC-M2-3 NMOS_OR1 l=1u w=2u
M4 NC-M4-0 NC-M4-1 NC-M4-2 NC-M4-3 NMOS_OR1 l=1u w=2u
M6 NC-M6-0 NC-M6-1 NC-M6-2 NC-M6-3 NMOS_OR1 l=1u w=2u

.ends
