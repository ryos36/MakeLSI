.title KiCad schematic
M15 Net-_M15-Pad1_ /Vin1 Net-_M15-Pad3_ /VDD PMOS l=1u w=2u
M16 Net-_M15-Pad1_ /Vin1 Net-_M16-Pad3_ /Vss NMOS l=1u w=2u
M17 Net-_M15-Pad3_ Net-_M15-Pad1_ /VDD /VDD PMOS l=1u w=2u
M18 Net-_M16-Pad3_ Net-_M15-Pad1_ /Vss /Vss NMOS l=1u w=2u
M19 Net-_M19-Pad1_ /Vin2 Net-_M15-Pad3_ /VDD PMOS l=1u w=2u
M20 Net-_M19-Pad1_ /Vin2 Net-_M16-Pad3_ /Vss NMOS l=1u w=2u
M21 /Vout Net-_M19-Pad1_ /VDD /VDD PMOS l=1u w=6u
M22 /Vout Net-_M19-Pad1_ /Vss /Vss NMOS l=1u w=2u
.end
